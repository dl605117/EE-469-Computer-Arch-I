module fetch (


)

endmodule
