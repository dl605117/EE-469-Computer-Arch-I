module mem (


)

endmodule
