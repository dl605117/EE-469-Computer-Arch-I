module write_back (


)

endmodule
