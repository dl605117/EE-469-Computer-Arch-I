module execute (


)

endmodule
