module decode_reg_r (


)

endmodule
